// Simple 2-input AND gate
module and_gate(input wire A, B, output wire Y);
  assign Y = A & B;
endmodule